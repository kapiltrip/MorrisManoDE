module 
    //does nothing 
endmodule 